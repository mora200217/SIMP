// Module for flex senssor reading adc via SPI 
module flex_sensor (
    input rst, 
    

    output decod 

);
    
endmodule