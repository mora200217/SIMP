module segment_display(
    input [6:0] value, // 7 bits -> 0 - 127
    
); 

// convert value into d c u 



endmodule